Vcc 1 0 0
GB 6 3 (2,5) 7.294236337m
Vd 7 4 0
HD 5 8 Vd 8.389800025k
R1 2 1 1.017479474k
R2 2 3 2.034385969k
R3 2 5 3.084568126k
R4 0 5 4.169099379k
R5 6 5 3.007681327k
R6 0 7 2.042113276k
R7 4 8 1.005870522k
C 6 8 1.035738228u
.op
.ic V(6)=8.523047 v(8)=1.776357e-15
.end
